.SUBCKT OPAMP vip vin 4 1 7
* vip vip 
* vin vin
* 4 vout
* 1 VDD
* 7 VSS

M1 6 vin 3 3 p08 W=6U L=1U 
M2 5 vip 3 3 p08 W=6U L=1U
M3 6 6 7 7 n08 W=7U L=1U  
M4 5 6 7 7 n08 W=7U L=1U 
M5 3 2 1 1 p08 W=11U L=1U 
M6 4 5 7 7 n08 W=44U L=1U 
M7 4 2 1 1 p08 W=34U L=1U 
M8 2 2 1 1 p08 W=11U L=1U
Cc 4 5 3p
IR 2 7 30u


.MODEL n08 NMOS VTO = 0.70 KP = 110U GAMMA = 0.4  LAMBDA = 0.04 
+ PHI = 0.7 MJ = 0.5 MJSW = 0.38 CGBO = 700P CGSO = 220P CGDO = 220P 
+ CJ = 770U CJSW = 380P LD = 0.016U TOX = 14N
.MODEL p08 PMOS VTO = -0.70 KP = 50U GAMMA = 0.57 LAMBDA = 0.05 
+ PHI = 0.8 MJ = 0.5 MJSW = 0.35 CGBO = 700P CGSO = 220P CGDO = 220P 
+ CJ = 560U CJSW = 350P LD = 0.014U TOX = 14N

.ENDS